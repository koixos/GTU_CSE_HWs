module cla_16bit (
	output [15:0] sum,
	output cout,
	input [15:0] ain,
	input [15:0] bin,
	input cin
);
	
	wire [15:0] prop;
	wire [15:0] gen;
	wire carry;
	
	cla_8bit cla1 (
		.sum(sum[7:0]),
		.cout(carry),
		.ain(ain[7:0]),
		.bin(bin[7:0]),
		.cin(cin)
	);
	
	cla_8bit cla2 (
		.sum(sum[15:8]),
		.cout(cout),
		.ain(ain[15:8]),
		.bin(bin[15:8]),
		.cin(carry)
	);
	
endmodule